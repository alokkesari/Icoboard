module not_module(input a, output out);
assign out=~a;
endmodule
